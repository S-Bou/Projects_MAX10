-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Mon Feb 15 19:13:40 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY P_3 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        MONO : IN STD_LOGIC := '0';
        EQUAL : IN STD_LOGIC := '0';
        OPERATE : OUT STD_LOGIC;
        ALARM : OUT STD_LOGIC
    );
END P_3;

ARCHITECTURE BEHAVIOR OF P_3 IS
    TYPE type_fstate IS (Q0,Q1,Q2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,MONO,EQUAL)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Q0;
            OPERATE <= '0';
            ALARM <= '0';
        ELSE
            OPERATE <= '0';
            ALARM <= '0';
            CASE fstate IS
                WHEN Q0 =>
                    IF ((NOT((MONO = '1')) AND (EQUAL = '1'))) THEN
                        reg_fstate <= Q1;
                    ELSIF ((NOT((MONO = '1')) AND NOT((EQUAL = '1')))) THEN
                        reg_fstate <= Q2;
                    ELSE
                        reg_fstate <= Q0;
                    END IF;

                    OPERATE <= '0';

                    ALARM <= '0';
                WHEN Q1 =>
                    IF (((MONO = '1') AND NOT((EQUAL = '1')))) THEN
                        reg_fstate <= Q0;
                    ELSIF ((NOT((MONO = '1')) AND NOT((EQUAL = '1')))) THEN
                        reg_fstate <= Q2;
                    ELSE
                        reg_fstate <= Q1;
                    END IF;

                    OPERATE <= '0';

                    ALARM <= '1';
                WHEN Q2 =>
                    IF (((NOT((MONO = '1')) AND (EQUAL = '1')) OR ((MONO = '1') AND (EQUAL = '1')))) THEN
                        reg_fstate <= Q0;
                    ELSE
                        reg_fstate <= Q2;
                    END IF;

                    OPERATE <= '1';

                    ALARM <= '0';
                WHEN OTHERS => 
                    OPERATE <= 'X';
                    ALARM <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
