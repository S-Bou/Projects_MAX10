library ieee; 
use ieee.std_logic_1164.all;
use work.mux4to1_package.all;

entity Step_Motor_Driver is

end Step_Motor_Driver;