-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Sun Feb 28 13:47:33 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        Pulse : IN STD_LOGIC := '0';
        Led_9 : OUT STD_LOGIC;
        Led_8 : OUT STD_LOGIC;
        Led_7 : OUT STD_LOGIC;
        Led_6 : OUT STD_LOGIC
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (Q0,Q1,Q2,Q3,Q4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Pulse)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Q0;
            Led_9 <= '0';
            Led_8 <= '0';
            Led_7 <= '0';
            Led_6 <= '0';
        ELSE
            Led_9 <= '0';
            Led_8 <= '0';
            Led_7 <= '0';
            Led_6 <= '0';
            CASE fstate IS
                WHEN Q0 =>
                    IF ((Pulse = '1')) THEN
                        reg_fstate <= Q1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Q0;
                    END IF;
                WHEN Q1 =>
                    IF ((Pulse = '1')) THEN
                        reg_fstate <= Q2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Q1;
                    END IF;

                    Led_9 <= '1';
                WHEN Q2 =>
                    IF ((Pulse = '1')) THEN
                        reg_fstate <= Q3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Q2;
                    END IF;

                    Led_8 <= '1';
                WHEN Q3 =>
                    IF ((Pulse = '1')) THEN
                        reg_fstate <= Q4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Q3;
                    END IF;

                    Led_7 <= '1';
                WHEN Q4 =>
                    IF ((Pulse = '1')) THEN
                        reg_fstate <= Q0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Q4;
                    END IF;

                    Led_6 <= '1';
                WHEN OTHERS => 
                    Led_9 <= 'X';
                    Led_8 <= 'X';
                    Led_7 <= 'X';
                    Led_6 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
